module Adder ();

endmodule // Adder

module Accumulator ();

endmodule // Accumulator

module Adder ();
  
endmodule // Adder
